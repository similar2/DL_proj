module jump(
    input en,
    input [7:0] i_num,
    input [1:0] func,
    input clk,
    input [7:0] feedbak_sig,//current state in the kitchen
    output [4:0] control_data //control when to do the movement i.e. get put etc
);



endmodule