`timescale 1ns/1ps

module TravelerOperateMachine(
    input button_left,      // get
    input button_center,    // move
    input button_right,     // put
    input switch_right_0,   // interact
    input switch_right_1,    // throw
    input output_ready,
    output reg [7:0] output_data
);
always@(*)
begin
end



endmodule