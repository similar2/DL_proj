`timescale 1ns/1ps

module ChangeTargetMachine(
    input button_up,
    input button_down,
    input output_ready,
    output reg [7:0] output_data
);

endmodule