`timescale 1ns/1ps

module ChangeGameState(
    input switch_left_0,
    input output_ready,
    output reg [7:0] output_data
);

endmodule